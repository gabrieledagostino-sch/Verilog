module XOR4(z,a);
    output     z;
    input [3:0]a;

    assign z = (~a[0] &  a[1] &  a[2] &  a[3]) | ( a[0] & ~a[1] &  a[2] &   a[3]) |
               ( a[0] &  a[1] & ~a[2] &  a[3]) | ( a[0] &  a[1] &  a[2] &  ~a[3]) |
               (~a[0] & ~a[1] & ~a[2] &  a[3]) | (~a[0] & ~a[1] &  a[2] &  ~a[3]) |
               (~a[0] &  a[1] & ~a[2] & ~a[3]) | ( a[0] & ~a[1] & ~a[2] &  ~a[3]) ;
endmodule